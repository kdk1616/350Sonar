`timescale 1ns / 1ps
/**
 * 
 * READ THIS DESCRIPTION:
 *
 * This is the Wrapper module that will serve as the header file combining your processor, 
 * RegFile and Memory elements together.
 *
 * This file will be used to generate the bitstream to upload to the FPGA.
 * We have provided a sibling file, Wrapper_tb.v so that you can test your processor's functionality.
 * 
 * We will be using our own separate Wrapper_tb.v to test your code. You are allowed to make changes to the Wrapper files 
 * for your own individual testing, but we expect your final processor.v and memory modules to work with the 
 * provided Wrapper interface.
 * 
 * Refer to Lab 5 documents for detailed instructions on how to interface 
 * with the memory elements. Each imem and dmem modules will take 12-bit 
 * addresses and will allow for storing of 32-bit values at each address. 
 * Each memory module should receive a single clock. At which edges, is 
 * purely a design choice (and thereby up to you). 
 * 
 * You must change line 36 to add the memory file of the test you created using the assembler
 * For example, you would add sample inside of the quotes on line 38 after assembling sample.s
 *
 **/

module FPGAWrapper (
    input CLK100MHZ, 
    input CPU_RESETN, 
    output[7:0] LED, 
    inout[15:0] PINS,
    output hSync, 		// H Sync Signal
	output vSync, 		// Veritcal Sync Signal
	output[3:0] VGA_R,  // Red Signal Bits
	output[3:0] VGA_G,  // Green Signal Bits
	output[3:0] VGA_B  // Blue Signal Bits
	);
	
	wire reset = ~CPU_RESETN;;

	wire rwe, mwe;
	wire[4:0] rd, rs1, rs2;
	wire[31:0] instAddr, instData, 
		rData, regA, regB,
		memAddr, memDataIn, memDataOut;


	wire CLK;
	tff clock_tff(CLK, 1'b1, CLK100MHZ, 1'b0);
	

	// ADD YOUR MEMORY FILE HERE
	localparam INSTR_FILE = "read_seq";
	
	// Main Processing Unit
	processor CPU(
		// .debug(debug),
		.clock(CLK), .reset(reset), 
								
		// ROM
		.address_imem(instAddr), .q_imem(instData),
									
		// Regfile
		.ctrl_writeEnable(rwe),     .ctrl_writeReg(rd),
		.ctrl_readRegA(rs1),     .ctrl_readRegB(rs2), 
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB),
									
		// RAM
		.wren(mwe), .address_dmem(memAddr), 
		.data(memDataIn), .q_dmem(memDataOut),
		
		.io_pins(PINS)); 
	
	assign LED[7:0] = memAddr;
	
	// Instruction Memory (ROM)
	ROM #(.MEMFILE({INSTR_FILE, ".mem"}))
	InstMem(.clk(CLK), 
		.addr(instAddr[11:0]), 
		.dataOut(instData));
	
	// Register File
	regfile RegisterFile(.clock(CLK), 
		.ctrl_writeEnable(rwe), .ctrl_reset(reset), 
		.ctrl_writeReg(rd),
		.ctrl_readRegA(rs1), .ctrl_readRegB(rs2), 
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB));
						

	// Processor Memory (RAM)
	RAM ProcMem(.clk(CLK), 
		.wEn(mwe), 
		.addr(memAddr[11:0]), 
		.dataIn(memDataIn), 
		.dataOut(memDataOut)
	);


	wire[18:0] vgaPixelAddr, cpuPixelAddr;
	wire vgaPixelOut, cpuPixelOut;
	wire cpuPixelIn;
	wire pixel_wEn = 1'b0;


	DPRAM #(
		.DEPTH(640*480), 		       // Set depth to contain every color		
		.DATA_WIDTH(1), 		       // Set data width according to the bits per color
		.ADDRESS_WIDTH(19)     // Set address width according to the color count
		)  // Memory initialization
	pixelRam(
		.clk(CLK), 	
		.wEn0(pixel_wEn),
		.wEn1(1'b0),	
		.addr0(cpuPixelAddr),
		.addr1(vgaPixelAddr),
		.dataIn0(cpuPixelIn),
		.dataIn1(1'b0),
		.dataOut0(cpuPixelOut),
		.dataOut0(vgaPixelOut)
	); 
	
	VGAController vga(     
	CLK100MHZ, 			// 100 MHz System Clock
	CPU_RESETN, 		// Reset Signal
	hSync, 		// H Sync Signal
	vSync, 		// Veritcal Sync Signal
	VGA_R,  // Red Signal Bits
	VGA_G,  // Green Signal Bits
	VGA_B,  // Blue Signal Bits
	pixelAddr,
	pixelOut
	);
		
endmodule